module keyboard(
    input[6:0] key,
    output pwm
);

endmodule