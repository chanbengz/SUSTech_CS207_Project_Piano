module learning(
	input clk,
    input [7:0] key,
	input [2:0] mode,
	input [1:0] song_num,
	output speaker,
	output reg [7:0] led,
	output reg [3:0] pitch
	);

endmodule