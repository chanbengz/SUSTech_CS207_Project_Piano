module sig_sel(
    input clk, rst_n,
    input [2:0] mode,
    input [1:0] song_num,
    input speaker1, speaker2, speaker3,
    input [7:0] led1, led2,
    output reg speaker,
    output [7:0] seg_en, [7:0] seg_out0, seg_out1,
    output reg led
    );

     reg [3:0] p0, p1, p2, p3, p4, p5, p6, p7;
     seg_display(.clk(clk),
                 .rst_n(rst_n),
                 .p0(p0),.p1(p1),.p2(p2),.p3(p3),.p4(p4),.p5(p5),.p6(p6),.p7(p7),
                 .seg_en(seg_en),.seg_out0(seg_out0), .seg_out1(seg_out1)
                 );

    always @(posedge clk) begin
        case(mode)
            3'b011: begin
                p7 <= 'hA;
                p6 <= {2'b00, song_num};
                {p5, p4, p3, p2, p1, p0} <= 'hDDDDDD;
                led <= led1;
                speaker <= speaker1;
            end
            3'b001: begin
                {p7, p6, p5, p4} <= 'hF4EE;
                {p3, p2, p1, p0} <= 'hDDDD;
                led <= 8'b0000_0000;
                speaker <= speaker2;
            end
            3'b111: begin
                led <= led2;
                speaker <= speaker3;
            end
            default: begin
                {p7, p6, p5, p4, p3} <= 'h5E660; // hello message
                {p2, p1, p0} <= 'hDDD;
                led <= 8'b0000_0000;
                speaker <= 0;
            end
        endcase
    end

endmodule