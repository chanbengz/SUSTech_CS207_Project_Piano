module sig_sel(
    input [2:0] mode,
    input sig1, sig2, sig3,
    output reg sig_out
    );

endmodule