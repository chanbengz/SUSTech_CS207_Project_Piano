module sig_sel(
    input [2:0] mode,
    input [1:0] song_num,
    input sig1, sig2, sig3,
    output reg sig_out,
    output reg [7:0] seg_en, seg_out0, seg_out1
    );

endmodule